module OR(output out1,  input in1, in2);
  or (out1, in1, in2);
endmodule
